//////////////////////////////////////////////////////////////////////////////////
// Test bench for Exercise #8 - Times Table using AXI interface
// Student Name: Ben Kaye
// Date: 2020-06-03
//
// Description: A testbench module to test Ex8 - Times Table using AXI4-Lite
// You need to write the whole file
//////////////////////////////////////////////////////////////////////////////////

//MIGHT HAVE TO CHANGE THE TIME SCALE
`timescale 1ns / 100ps

module test();
	//MAY NEED TO MOD
	parameter CLK_PRD = 4;
	
	reg clk, rst, read, err, t;
	reg [2:0] a, b, d;
	wire [5:0] result; 

	initial begin
		rst <= 0;
		err <= 0;
		clk <= 0;
		read <= 0;
		err <= 0;
		a <= 3'd3;
		b <= 3'd7;
		d <= 3'd3;
		forever #(CLK_PRD/2) clk = ~clk;
	end

    always  @(posedge clk) begin
            
            err <= (result != a*b && d==3'd3)  ? 1 : err;
            
            a <= (d==3'd3) ? {$random} % 8 : a;
            b <= (d==3'd3) ? {$random} % 8 : b;
            read <= d[1];
            
            
		
            d[2:1]<=d[1:0];
            d[0] <= d[2];
            
        
    end
    
	initial begin
		#400 begin 
			if (err) $display("Error encountered.");
			else $display("No error detected.");
			$finish; 
		end
	end
    
	axi_multiplier mplier(
		.a(a),
		.b(b),
		.clk(clk),
		.rst(rst),
		.read(read),
		.result(result)
	);
endmodule
